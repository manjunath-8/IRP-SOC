--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%% 
--%%                      Centre for Development of Advanced Computing                            %%
--%%                           Vellayambalam, Thiruvananthapuram.                                 %%
--%%==============================================================================================%%
--%% This confidential and proprietary software may be used only as authorised by a licensing     %%
--%% agreement from Centre for Development of Advanced Computing, India (C-DAC).In the event of   %%
--%% publication, the following notice is applicable:                                             %%
--%% Copyright (c) 2024 C-DAC                                                                     %%
--%% ALL RIGHTS RESERVED                                                                          %%
--%% The entire notice above must be reproduced on all authorised copies.                         %%
--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
--%% Project  Name    : Development of 32-bit RISC-V processor (RV32IM)                           %%
--%% Project Code     : HDG083D                                                                   %%
--%% File Name        : ROM_32KB_TOP.vhdl                                                         %%
--%% Title            :                                                                           %%
--%% Author           : vega@cdac.in                                                              %%               
--%% Description      : Top file that sends and receives the read signals from ROM controller     %%
---%% Version          : 00                                                                       %%
--%%%%%%%%%%%%%%%%%%%% Modification / Updation  History %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

----%% Date----------By---------------Version----Change Description-------------------------------%%
----%%                                                                                            %%
----%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ROM_THEJAS32 is
	Port (	
			clk		: IN STD_LOGIC;
	        rst_n   : IN STD_LOGIC;
			ena     : IN STD_LOGIC;
       		addra   : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
       		douta   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
       		enb     : IN STD_LOGIC;
       		addrb   : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
       		doutb   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)

		 );
end ROM_THEJAS32;

architecture ROM_THEJAS32_a of ROM_THEJAS32 is

	type rom_type is array(0 to 1972) of STD_LOGIC_VECTOR(31 DOWNTO 0);
	constant CDAC_rom	:	rom_type:=(
"00000000000000000000000010010011",                                                                                                
"00000000000000000000000100010011",                                                                                                
"00000000000000000000000110010011",                                                                                                
"00000000000000000000001000010011",                                                                                                
"00000000000000000000001010010011",                                                                                                
"00000000000000000000001100010011",                                                                                                
"00000000000000000000001110010011",                                                                                                
"00000000000000000000010000010011",                                                                                                
"00000000000000000000010010010011",                                                                                                
"00000000000000000000010100010011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000000000000011000010011",                                                                                                
"00000000000000000000011010010011",                                                                                                
"00000000000000000000011100010011",                                                                                                
"00000000000000000000011110010011",                                                                                                
"00000000000000000000100000010011",                                                                                                
"00000000000000000000100010010011",                                                                                                
"00000000000000000000100100010011",                                                                                                
"00000000000000000000100110010011",                                                                                                
"00000000000000000000101000010011",                                                                                                
"00000000000000000000101010010011",                                                                                                
"00000000000000000000101100010011",                                                                                                
"00000000000000000000101110010011",                                                                                                
"00000000000000000000110000010011",                                                                                                
"00000000000000000000110010010011",                                                                                                
"00000000000000000000110100010011",                                                                                                
"00000000000000000000110110010011",                                                                                                
"00000000000000000000111000010011",                                                                                                
"00000000000000000000111010010011",                                                                                                
"00000000000000000000111100010011",                                                                                                
"00000000000000000000111110010011",                                                                                                
"00000000000100000000001010010011",                                                                                                
"00000001111100101001001010010011",                                                                                                
"00000000000000101100010001100011",                                                                                                
"00000000000000000000000001101111",                                                                                                
"00000000000000000000001010010111",                                                                                                
"00001000000000101000001010010011",                                                                                                
"00110000010100101001000001110011",                                                                                                
"00000000001000101111000110010111",                                                                                                
"11111000000000011000000110010011",                                                                                                
"10101110100100011000001000010011",                                                                                                
"11111100000000100111001000010011",                                                                                                
"00000000000100000000011010010011",                                                                                                
"10000000100000011000010110010011",                                                                                                
"00000000110101011010000000100011",                                                                                                
"11110001010000000010010101110011",                                                                                                
"00000010000001010000111001100011",                                                                                                
"00000000000100000000010110010011",                                                                                                
"00000000101101010111000001100011",                                                                                                
"00000000000100000000011010010011",                                                                                                
"10000000100000011000010110010011",                                                                                                
"00000000000001011010011000000011",                                                                                                
"11111110110101100000110011100011",                                                                                                
"11110001010000000010010101110011",                                                                                                
"11000000000000000000010110110111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000001000000001111",                                                                                                
"00001111111100000000000000001111",                                                                                                
"10000000000000000000011000110111",                                                                                                
"00000000000001100000000001100111",                                                                                                
"00000000110001010001011000010011",                                                                                                
"00000000110000100000001000110011",                                                                                                
"00000000000101010000000100010011",                                                                                                
"00000000110000010001000100010011",                                                                                                
"00000000010000010000000100110011",                                                                                                
"00101101100000000000000001101111",                                                                                                
"11101111000000010000000100010011",                                                                                                
"00000000000100010010001000100011",                                                                                                
"00000000001000010010010000100011",                                                                                                
"00000000001100010010011000100011",                                                                                                
"00000000010000010010100000100011",                                                                                                
"00000000010100010010101000100011",                                                                                                
"00000000011000010010110000100011",                                                                                                
"00000000011100010010111000100011",                                                                                                
"00000010100000010010000000100011",                                                                                                
"00000010100100010010001000100011",                                                                                                
"00000010101000010010010000100011",                                                                                                
"00000010101100010010011000100011",                                                                                                
"00000010110000010010100000100011",                                                                                                
"00000010110100010010101000100011",                                                                                                
"00000010111000010010110000100011",                                                                                                
"00000010111100010010111000100011",                                                                                                
"00000101000000010010000000100011",                                                                                                
"00000101000100010010001000100011",                                                                                                
"00000101001000010010010000100011",                                                                                                
"00000101001100010010011000100011",                                                                                                
"00000101010000010010100000100011",                                                                                                
"00000101010100010010101000100011",                                                                                                
"00000101011000010010110000100011",                                                                                                
"00000101011100010010111000100011",                                                                                                
"00000111100000010010000000100011",                                                                                                
"00000111100100010010001000100011",                                                                                                
"00000111101000010010010000100011",                                                                                                
"00000111101100010010011000100011",                                                                                                
"00000111110000010010100000100011",                                                                                                
"00000111110100010010101000100011",                                                                                                
"00000111111000010010110000100011",                                                                                                
"00000111111100010010111000100011",                                                                                                
"00110100001000000010010101110011",                                                                                                
"00110100000100000010010111110011",                                                                                                
"00000000000000010000011000010011",                                                                                                
"00001001100000000000000011101111",                                                                                                
"00110100000101010001000001110011",                                                                                                
"00000000000000000010001010110111",                                                                                                
"10000000000000101000001010010011",                                                                                                
"00110000000000101010000001110011",                                                                                                
"00000000010000010010000010000011",                                                                                                
"00000000100000010010000100000011",                                                                                                
"00000000110000010010000110000011",                                                                                                
"00000001000000010010001000000011",                                                                                                
"00000001010000010010001010000011",                                                                                                
"00000001100000010010001100000011",                                                                                                
"00000001110000010010001110000011",                                                                                                
"00000010000000010010010000000011",                                                                                                
"00000010010000010010010010000011",                                                                                                
"00000010100000010010010100000011",                                                                                                
"00000010110000010010010110000011",                                                                                                
"00000011000000010010011000000011",                                                                                                
"00000011010000010010011010000011",                                                                                                
"00000011100000010010011100000011",                                                                                                
"00000011110000010010011110000011",                                                                                                
"00000100000000010010100000000011",                                                                                                
"00000100010000010010100010000011",                                                                                                
"00000100100000010010100100000011",                                                                                                
"00000100110000010010100110000011",                                                                                                
"00000101000000010010101000000011",                                                                                                
"00000101010000010010101010000011",                                                                                                
"00000101100000010010101100000011",                                                                                                
"00000101110000010010101110000011",                                                                                                
"00000110000000010010110000000011",                                                                                                
"00000110010000010010110010000011",                                                                                                
"00000110100000010010110100000011",                                                                                                
"00000110110000010010110110000011",                                                                                                
"00000111000000010010111000000011",                                                                                                
"00000111010000010010111010000011",                                                                                                
"00000111100000010010111100000011",                                                                                                
"00000111110000010010111110000011",                                                                                                
"00010001000000010000000100010011",                                                                                                
"00110000001000000000000001110011",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110101101000010010000100011",                                                                                                
"11111110110001000010001000100011",                                                                                                
"00000000000000000001010100010111",                                                                                                
"01110010000001010000010100010011",                                                                                                
"01000111000000000000000011101111",                                                                                                
"00000000000000000000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111111000000010000000100010011",                                                                                                
"00000000000100010010011000100011",                                                                                                
"00000000100000010010010000100011",                                                                                                
"00000001000000010000010000010011",                                                                                                
"00000000000000000001010100010111",                                                                                                
"01101111100001010000010100010011",                                                                                                
"01000011110000000000000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000110000010010000010000011",                                                                                                
"00000000100000010010010000000011",                                                                                                
"00000001000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"00000000000000000001010100010111",                                                                                                
"01101100110001010000010100010011",                                                                                                
"01000000100000000000000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000100000010010111000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110101101000010010000100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"11111110000001111001111011100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110101101000010010000100011",                                                                                                
"00000000000000000001010100010111",                                                                                                
"01100110100001010000010100010011",                                                                                                
"11110111100111111111000011101111",                                                                                                
"11111111111100000000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"01001011000001111010011110000011",                                                                                                
"00000000010001111000011110110011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"01001010010001111010011110000011",                                                                                                
"00000000010001111000011110110011",                                                                                                
"01000000111101110000011110110011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"00000000000000100000011110010011",                                                                                                
"11111110110001000010011000000011",                                                                                                
"10101010101000011000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00001010010000000000000011101111",                                                                                                
"00000000001000101110011110010111",                                                                                                
"01001000000001111010011110000011",                                                                                                
"00000000010001111000011110110011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"01000110100001111010011110000011",                                                                                                
"00000000010001111000011110110011",                                                                                                
"01000000111101110000011110110011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"00000000000000100000011100010011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110100001000010011000000011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00010100000000000000000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11110100110111111111000011101111",                                                                                                
"11111101100001000010010110000011",                                                                                                
"11111101110001000010010100000011",                                                                                                
"11101101000111111111000011101111",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000000000000010100010011",                                                                                                
"00111100000000000001000011101111",                                                                                                
"11111110101001000010011000100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111100110001000010101000100011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"00000000111101110110011100110011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000111101110110011110110011",                                                                                                
"00000000001101111111011110010011",                                                                                                
"00000100000001111001100001100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"00000010010000000000000001101111",                                                                                                
"11111110110001000010011100000011",                                                                                                
"00000000010001110000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000010001111000011010010011",                                                                                                
"11111110110101000010010000100011",                                                                                                
"00000000000001110010011100000011",                                                                                                
"00000000111001111010000000100011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110100001000010011100000011",                                                                                                
"11111100111101110110100011100011",                                                                                                
"00000100110000000000000001101111",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111110111101000010001000100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"11111110111101000010000000100011",                                                                                                
"00000010010000000000000001101111",                                                                                                
"11111110010001000010011100000011",                                                                                                
"00000000000101110000011110010011",                                                                                                
"11111110111101000010001000100011",                                                                                                
"11111110000001000010011110000011",                                                                                                
"00000000000101111000011010010011",                                                                                                
"11111110110101000010000000100011",                                                                                                
"00000000000001110100011100000011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110000001000010011100000011",                                                                                                
"11111100111101110110100011100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111100110001000010101000100011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000111101110110011110110011",                                                                                                
"00000000001101111111011110010011",                                                                                                
"00000110000001111001100001100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"00001111111101111111011110010011",                                                                                                
"11111110111101000010001000100011",                                                                                                
"11111110010001000010011110000011",                                                                                                
"00000000100001111001011110010011",                                                                                                
"11111110010001000010011100000011",                                                                                                
"00000000111101110110011110110011",                                                                                                
"11111110111101000010001000100011",                                                                                                
"11111110010001000010011110000011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"11111110010001000010011100000011",                                                                                                
"00000000111101110110011110110011",                                                                                                
"11111110111101000010001000100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"00000001100000000000000001101111",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000010001111000011100010011",                                                                                                
"11111110111001000010011000100011",                                                                                                
"11111110010001000010011100000011",                                                                                                
"00000000111001111010000000100011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110110001000010011100000011",                                                                                                
"11111100111101110110111011100011",                                                                                                
"00000011110000000000000001101111",                                                                                                
"11111101110001000010011110000011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"00000001110000000000000001101111",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000000101111000011100010011",                                                                                                
"11111110111001000010010000100011",                                                                                                
"11111101100001000010011100000011",                                                                                                
"00001111111101110111011100010011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110100001000010011100000011",                                                                                                
"11111100111101110110110011100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000100000010010111000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00001000001100000000011100010011",                                                                                                
"00000000111001111010011000100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000111001111010000000100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000000000001111010001000100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000000001100000000011100010011",                                                                                                
"00000000111001111010011000100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000000000001111010001000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100111101000000111110100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000111001111010000000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000001010001111010011110000011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000010000001111111011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000010000000000000011110010011",                                                                                                
"11111100111101110001110011100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"00000010000000000000000001101111",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110111010111111111000011101111",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"11111100000001111001111011100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000100000010010111000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000001010001111010011110000011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000101111111011110010011",                                                                                                
"11111110000001111000001011100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000000000001111010011110000011",                                                                                                
"11111110111101000000011100100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"11111110111001000100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000001110000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111110000001000001011100100011",                                                                                                
"11111110000001000010010000100011",                                                                                                
"00001010110000000000000001101111",                                                                                                
"11111101110001000010011100000011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000100001111001011110010011",                                                                                                
"00000001000001111001011100010011",                                                                                                
"01000001000001110101011100010011",                                                                                                
"11111110111001000001011110000011",                                                                                                
"00000000111101110100011110110011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"00000000100000000000011110010011",                                                                                                
"11111110111101000000001110100011",                                                                                                
"00000101110000000000000001101111",                                                                                                
"11111110111001000001011110000011",                                                                                                
"00000010000001111101111001100011",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000000101111001011110010011",                                                                                                
"00000001000001111001011100010011",                                                                                                
"01000001000001110101011100010011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"00000011100001111000011110010011",                                                                                                
"00000000000001111101011110000011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"00000000111101110100011110110011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"00000001000000000000000001101111",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000000101111001011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"11111110011101000100011110000011",                                                                                                
"11111111111101111000011110010011",                                                                                                
"11111110111101000000001110100011",                                                                                                
"11111110011101000100011110000011",                                                                                                
"11111010000001111001001011100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111110100001000010011100000011",                                                                                                
"11110100111101110110100011100011",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000100000010010111000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110000001000010010000100011",                                                                                                
"00001010110000000000000001101111",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"00000001000001111101011110010011",                                                                                                
"00000000100001111001011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"00000000100000000000011110010011",                                                                                                
"11111110111101000000001110100011",                                                                                                
"00000101110000000000000001101111",                                                                                                
"11111110111001000001011110000011",                                                                                                
"00000010000001111101111001100011",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000000101111001011110010011",                                                                                                
"00000001000001111001011100010011",                                                                                                
"01000001000001110101011100010011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"11110111100001111000011110010011",                                                                                                
"00000000000001111101011110000011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"00000000111101110100011110110011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"00000001000000000000000001101111",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000000101111001011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"11111110011101000100011110000011",                                                                                                
"11111111111101111000011110010011",                                                                                                
"11111110111101000000001110100011",                                                                                                
"11111110011101000100011110000011",                                                                                                
"11111010000001111001001011100011",                                                                                                
"00000000001000101110011100010111",                                                                                                
"11110100100001110000011100010011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000000101111001011110010011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110111001000101011100000011",                                                                                                
"00000000111001111001000000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111110100001000010011100000011",                                                                                                
"00001111111100000000011110010011",                                                                                                
"11110100111001111111100011100011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"11101111100001111000011110010011",                                                                                                
"00000000000100000000011100010011",                                                                                                
"00000000111001111010000000100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111100110001000010101000100011",                                                                                                
"11111100111101000001111100100011",                                                                                                
"11111101111001000101011110000011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"11101011000001111000011110010011",                                                                                                
"00000000000001111010011110000011",                                                                                                
"00000000000001111001010001100011",                                                                                                
"11101110000111111111000011101111",                                                                                                
"11111110000001000000011010100011",                                                                                                
"00000111110000000000000001101111",                                                                                                
"11111110110101000100011110000011",                                                                                                
"11111101100001000010011100000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000100001111101011110010011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"00000001000001111101011110010011",                                                                                                
"00000000111101110100011110110011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"00000000001000101110011100010111",                                                                                                
"11101000010001110000011100010011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000000101111001011110010011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"00000000000001111101011110000011",                                                                                                
"00000001000001111001011100010011",                                                                                                
"01000001000001110101011100010011",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000100001111001011110010011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"00000000111101110100011110110011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"01000001000001111101011110010011",                                                                                                
"11111110111101000001011100100011",                                                                                                
"11111110110101000100011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000000011010100011",                                                                                                
"11111110110101000100011110000011",                                                                                                
"11111101010001000010011100000011",                                                                                                
"11111000111001111110000011100011",                                                                                                
"11111110111001000101011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110101101000010010000100011",                                                                                                
"00000000000001100000011110010011",                                                                                                
"11111110111101000001001100100011",                                                                                                
"11111110011001000101011110000011",                                                                                                
"11111110100001000010011000000011",                                                                                                
"11111110110001000010010110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11101111000111111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100111101000000111110100011",                                                                                                
"11111110000001000000011110100011",                                                                                                
"11111110000001000010010000100011",                                                                                                
"11111101111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"00000011000000000000011110010011",                                                                                                
"00000000111101110010010000100011",                                                                                                
"11111110000001000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111111111111111110011110110111",                                                                                                
"00011111111101111000011110010011",                                                                                                
"00000000111101110111011110110011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"11101111111101111111011110010011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"11110011111101111111011110010011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"00000011000001111110011110010011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"11111111011101111111011110010011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"11111111101101111111011110010011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"11111111110001111111011110010011",                                                                                                
"11111110111101000001001000100011",                                                                                                
"11111101111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111110010001000101011110000011",                                                                                                
"00000000111101110001000000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100111101000000111110100011",                                                                                                
"11111110000001000000011110100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"11111101111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000010001111010011110000011",                                                                                                
"00000100000001111111011110010011",                                                                                                
"11111100000001111000000011100011",                                                                                                
"11111101111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000001000001111010011110000011",                                                                                                
"11111110111101000001011000100011",                                                                                                
"11111110110001000101011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"00000000000001011000011100010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00000000000001110000011110010011",                                                                                                
"11111110111101000001011000100011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00001010100000000000000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000010001111010011110000011",                                                                                                
"00001000000001111111011110010011",                                                                                                
"11111100000001111000000011100011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111110110001000101011110000011",                                                                                                
"00000000111101110010011000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000100000010010111000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000010001111010011110000011",                                                                                                
"00000001000001111111011110010011",                                                                                                
"11111100000001111001000011100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000100000010010111000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"00000000000001011000011100010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00000000000001110000011110010011",                                                                                                
"11111110111101000000011100100011",                                                                                                
"11111110111001000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00001000111101110001110001100011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000000001111101011110000011",                                                                                                
"00000001000001111001011100010011",                                                                                                
"00000001000001110101011100010011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011010000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101101001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011010000011",                                                                                                
"00000000000101101111011010010011",                                                                                                
"00000000100001101001011010010011",                                                                                                
"00000000110101111000011110110011",                                                                                                
"00000000000001111000011010010011",                                                                                                
"00010000000001110110011110010011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"00000001000001111101011110010011",                                                                                                
"00000000111101101001000000100011",                                                                                                
"00001001010000000000000001101111",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000101110111011100010011",                                                                                                
"00000000100001110001011100010011",                                                                                                
"00000000111001111000011110110011",                                                                                                
"00000000000001111101011110000011",                                                                                                
"00000001000001111001011100010011",                                                                                                
"00000001000001110101011100010011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"11111110111101000100011010000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101101001100001100011",                                                                                                
"00010000000000000000011110110111",                                                                                                
"01100000000001111000011110010011",                                                                                                
"00000000110000000000000001101111",                                                                                                
"00010000001000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"11111110111101000100011010000011",                                                                                                
"00000000000101101111011010010011",                                                                                                
"00000000100001101001011010010011",                                                                                                
"00000000110101111000011110110011",                                                                                                
"00000000000001111000011010010011",                                                                                                
"11101111111101110111011110010011",                                                                                                
"00000001000001111001011110010011",                                                                                                
"00000001000001111101011110010011",                                                                                                
"00000000111101101001000000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111100000000010000000100010011",                                                                                                
"00000010000100010010111000100011",                                                                                                
"00000010100000010010110000100011",                                                                                                
"00000100000000010000010000010011",                                                                                                
"11111100101001000010011000100011",                                                                                                
"11111110000001000010011000100011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111100000001000010110000100011",                                                                                                
"11111110000001000010001000100011",                                                                                                
"11111100000001000000111110100011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"10010000110001111000011110010011",                                                                                                
"00000000000001111010000000100011",                                                                                                
"00000000001000101110011110010111",                                                                                                
"10010000010001111000011110010011",                                                                                                
"00000000000000000001011100110111",                                                                                                
"00000010000101110000011100010011",                                                                                                
"00000000111001111001000000100011",                                                                                                
"00000101100000000000000001101111",                                                                                                
"00000100001100000000010100010011",                                                                                                
"11110010100011111111000011101111",                                                                                                
"11111110000001000010000000100011",                                                                                                
"00000011100000000000000001101111",                                                                                                
"00010000000000000000011110110111",                                                                                                
"00010000000001111000011110010011",                                                                                                
"00000001010001111010011110000011",                                                                                                
"11111100111101000000101110100011",                                                                                                
"11111101011101000100011110000011",                                                                                                
"00000000000101111111011110010011",                                                                                                
"00000000000001111000100001100011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"11111100111101000000111110100011",                                                                                                
"00000010000000000000000001101111",                                                                                                
"11111110000001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010000000100011",                                                                                                
"11111110000001000010011100000011",                                                                                                
"00000000000011110100011110110111",                                                                                                
"00100011111101111000011110010011",                                                                                                
"11111100111001111111000011100011",                                                                                                
"11111101111101000100011110000011",                                                                                                
"11111010000001111000010011100011",                                                                                                
"11111001000011111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"10100001110000011000011110010011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"10100001110000011000011110010011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000110111101110001001001100011",                                                                                                
"10100001110000011000010100010011",                                                                                                
"00010111110000000000000011101111",                                                                                                
"11111100110001000010011010000011",                                                                                                
"11111110110001000010011000000011",                                                                                                
"11111110100001000010010110000011",                                                                                                
"10100001110000011000010100010011",                                                                                                
"00001000010000000000000011101111",                                                                                                
"11111100101001000010110000100011",                                                                                                
"11111101100001000010011100000011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"11111010111101110000101011100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111110010001000010011110000011",                                                                                                
"00001000000001111000011110010011",                                                                                                
"11111110111101000010001000100011",                                                                                                
"11111110100001000010011100000011",                                                                                                
"00001111111100000000011110010011",                                                                                                
"11111000111001111111010011100011",                                                                                                
"11111110000001000010010000100011",                                                                                                
"11111000000111111111000001101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"10100001110000011000011110010011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"00000000010000000000011110010011",                                                                                                
"00000000111101110001101001100011",                                                                                                
"00000000011000000000010100010011",                                                                                                
"11100011010011111111000011101111",                                                                                                
"11111110010001000010011110000011",                                                                                                
"00000000100000000000000001101111",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000011110000010010000010000011",                                                                                                
"00000011100000010010010000000011",                                                                                                
"00000100000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111100110001000010101000100011",                                                                                                
"11111100110101000010100000100011",                                                                                                
"11111101100001000010010110000011",                                                                                                
"11111101110001000010010100000011",                                                                                                
"00011010000000000000000011101111",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110110001000010011100000011",                                                                                                
"11111111111100000000011110010011",                                                                                                
"00000110111101110000100001100011",                                                                                                
"11111110110001000010011100000011",                                                                                                
"11111111111000000000011110010011",                                                                                                
"00000110111101110000111001100011",                                                                                                
"11111110110001000010011100000011",                                                                                                
"11111111111000000000011110010011",                                                                                                
"00000110111001111110111001100011",                                                                                                
"11111110110001000010011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110000101001100011",                                                                                                
"11111110110001000010011100000011",                                                                                                
"11111111110100000000011110010011",                                                                                                
"00000100111101110000011001100011",                                                                                                
"00000110000000000000000001101111",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000001101111000011010010011",                                                                                                
"11111101010001000010011100000011",                                                                                                
"11111101000001000010011110000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"00000000000001111000010110010011",                                                                                                
"00000000000001101000010100010011",                                                                                                
"00001100110000000000000011101111",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00001000000001111000011110010011",                                                                                                
"11111100111101000010101000100011",                                                                                                
"00000000011000000000010100010011",                                                                                                
"11010111000011111111000011101111",                                                                                                
"00000010100000000000000001101111",                                                                                                
"00000001010100000000010100010011",                                                                                                
"11010110010011111111000011101111",                                                                                                
"00000001110000000000000001101111",                                                                                                
"00000001100000000000010100010011",                                                                                                
"11010101100011111111000011101111",                                                                                                
"00000001000000000000000001101111",                                                                                                
"00000000011000000000010100010011",                                                                                                
"11010100110011111111000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00000011010000000000000001101111",                                                                                                
"11011100110011111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"11111101110001000010011100000011",                                                                                                
"00000000111101110000011110110011",                                                                                                
"11111110100001000010011100000011",                                                                                                
"00001111111101110111011100010011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00001000010000000000011110010011",                                                                                                
"11111100111001111111010011100011",                                                                                                
"00000000000000000000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010100000010010011000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110000001000000010110100011",                                                                                                
"00000011100000000000000001101111",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111100111101000010111000100011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110101101000100011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000000010110100011",                                                                                                
"11111110101101000000011110000011",                                                                                                
"11111100000001111101010011100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111110000001000010011000100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"00000110111001111001010001100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000001001111000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000111101110000011100110011",                                                                                                
"00001111111100000000011110010011",                                                                                                
"00000010111101110001110001100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000001101111000011110010011",                                                                                                
"00001000001000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11001111000011111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000001111001011001100011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000011110000000000000001101111",                                                                                                
"11111111111100000000011110010011",                                                                                                
"00000011010000000000000001101111",                                                                                                
"11111111111100000000011110010011",                                                                                                
"00000010110000000000000001101111",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000011100010011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111111111101111000011110010011",                                                                                                
"00000000111101110001011001100011",                                                                                                
"11111111111000000000011110010011",                                                                                                
"00000000100000000000000001101111",                                                                                                
"11111111110100000000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100111101000000111110100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"11111101111101000100011100000011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110101010011111111000011101111",                                                                                                
"00001001111100000000011000010011",                                                                                                
"00000000001100000000010110010011",                                                                                                
"10101010010000011000010100010011",                                                                                                
"00100111000000000000000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01100111010001010000010100010011",                                                                                                
"10111001000011111111000011101111",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"00000001111100000000011110010011",                                                                                                
"00000010111101110001101001100011",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000000101111100011100000011",                                                                                                
"00001000011000000000011110010011",                                                                                                
"00000010111101110001001001100011",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000001001111100011100000011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"00000000111101110001101001100011",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01100100110001010000010100010011",                                                                                                
"10110101010011111111000011101111",                                                                                                
"00000101000000000000000001101111",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"00001011111100000000011110010011",                                                                                                
"00000010111101110001101001100011",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000000101111100011100000011",                                                                                                
"00000010010100000000011110010011",                                                                                                
"00000010111101110001001001100011",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000001001111100011100000011",                                                                                                
"00001000110100000000011110010011",                                                                                                
"00000000111101110001101001100011",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01100001100001010000010100010011",                                                                                                
"10110001010011111111000011101111",                                                                                                
"00000001000000000000000001101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01100001010001010000010100010011",                                                                                                
"10110000010011111111000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01100001010001010000010100010011",                                                                                                
"10101111100011111111000011101111",                                                                                                
"10101010010000011000011110010011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"00001011111100000000011110010011",                                                                                                
"00000100111101110001010001100011",                                                                                                
"11111000000000000000011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"10101010100000011000011110010011",                                                                                                
"00000101000000000000011100010011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"00000000000100000000010110010011",                                                                                                
"10101010100000011000010100010011",                                                                                                
"00101000000000000000000011101111",                                                                                                
"10101010100000011000011110010011",                                                                                                
"00000000000100000000011100010011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"10101010100000011000011110010011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000111001111000000010100011",                                                                                                
"00000000001000000000010110010011",                                                                                                
"10101010100000011000010100010011",                                                                                                
"00100101110000000000000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11111100101101000010110000100011",                                                                                                
"11111100110001000010101000100011",                                                                                                
"00000000001100000000011110010011",                                                                                                
"11111110111101000000011000100011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000001000001111101011110010011",                                                                                                
"00001111111101111111011110010011",                                                                                                
"11111110111101000000011010100011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00000000100001111101011110010011",                                                                                                
"00001111111101111111011110010011",                                                                                                
"11111110111101000000011100100011",                                                                                                
"11111101010001000010011110000011",                                                                                                
"00001111111101111111011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01010110100001010000010100010011",                                                                                                
"10100011010011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"10000111000111111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000100000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"10001100100111111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"11111110110001000100011100000011",                                                                                                
"00000000000001110000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110111000011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"11111110110101000100011100000011",                                                                                                
"00000000000001110000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110101100011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"11111110111001000100011100000011",                                                                                                
"00000000000001110000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110100000011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"11111110111101000100011100000011",                                                                                                
"00000000000001110000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110010100011111111000011101111",                                                                                                
"00000101000000000000000001101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110001000011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11100100110011111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"00001111111101111111011100010011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111100111101000010111000100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111111111101111000011110010011",                                                                                                
"11111100111101000010110000100011",                                                                                                
"11111101100001000010011110000011",                                                                                                
"11111010000001111001100011100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11111111110011111111000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110101101000010010000100011",                                                                                                
"00000000000001100000011110010011",                                                                                                
"11111110111101000000001110100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110100110011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000100000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11111010010011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"11111110011101000100011100000011",                                                                                                
"00000001000001110001011100010011",                                                                                                
"00000001000001110101011100010011",                                                                                                
"00000000000001110000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11100100010011111111000011101111",                                                                                                
"00000101000000000000000001101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11100010110011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11010110100011111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"00001111111101111111011100010011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000111001111000000000100011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"11111111111101111000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"11111010000001111001100011100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11110001100011111111000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"11111110101001000010011000100011",                                                                                                
"11111110101101000010010000100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11100111000011111111000011101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000100000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11101100100011111111000011101111",                                                                                                
"00000011100000000000000001101111",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011100000011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000001111000010110010011",                                                                                                
"00000000000001110000010100010011",                                                                                                
"11010110100011111111000011101111",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"11111111111101111000011110010011",                                                                                                
"11111110111101000010010000100011",                                                                                                
"11111110100001000010011110000011",                                                                                                
"11111100000001111001010011100011",                                                                                                
"10000000011000011000011110010011",                                                                                                
"00000000000001111100011110000011",                                                                                                
"00000000000000000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11100111010011111111000011101111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111110000000010000000100010011",                                                                                                
"00000000000100010010111000100011",                                                                                                
"00000000100000010010110000100011",                                                                                                
"00000010000000010000010000010011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"11111110111101000000011110100011",                                                                                                
"00000001100000000000000001101111",                                                                                                
"11111110111101000000011110010011",                                                                                                
"00000000010100000000011000010011",                                                                                                
"00000000000100000000010110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"11100100110111111111000011101111",                                                                                                
"11111110111101000100011110000011",                                                                                                
"00000000000101111111011110010011",                                                                                                
"11111110000001111001001011100011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000001110000010010000010000011",                                                                                                
"00000001100000010010010000000011",                                                                                                
"00000010000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111101000000010000000100010011",                                                                                                
"00000010000100010010011000100011",                                                                                                
"00000010100000010010010000100011",                                                                                                
"00000011000000010000010000010011",                                                                                                
"11111100101001000010111000100011",                                                                                                
"11110001010000000010010101110011",                                                                                                
"11111101110001000010011110000011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00000000000000000001000000001111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000000000000000000000000010011",                                                                                                
"10000000100000011000011110010011",                                                                                                
"00000000000001111010000000100011",                                                                                                
"00001111111100000000000000001111",                                                                                                
"00000000000000000001000000001111",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000001111000000011100111",                                                                                                
"00000000000000000000000000010011",                                                                                                
"00000010110000010010000010000011",                                                                                                
"00000010100000010010010000000011",                                                                                                
"00000011000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"11111100000000010000000100010011",                                                                                                
"00000010000100010010111000100011",                                                                                                
"00000010100000010010110000100011",                                                                                                
"00000100000000010000010000010011",                                                                                                
"10000000100000011000011110010011",                                                                                                
"00000000000100000000011100010011",                                                                                                
"00000000111001111010000000100011",                                                                                                
"11111110000001000010010000100011",                                                                                                
"11111110000001000010001000100011",                                                                                                
"11111110000001000010000000100011",                                                                                                
"00000000001000000000011110110111",                                                                                                
"11111100111101000010111000100011",                                                                                                
"11111100000001000000110110100011",                                                                                                
"00000000000100000000011110010011",                                                                                                
"11111100111101000010101000100011",                                                                                                
"00000000001000000000011110110111",                                                                                                
"11111100111101000010100000100011",                                                                                                
"00000001010100000000010100010011",                                                                                                
"11011101010111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00100000100001010000010100010011",                                                                                                
"11101010000111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00100000010001010000010100010011",                                                                                                
"11101001010111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00100100110001010000010100010011",                                                                                                
"11101000100111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00101001010001010000010100010011",                                                                                                
"11100111110111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00011110000001010000010100010011",                                                                                                
"11100111000111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00101101000001010000010100010011",                                                                                                
"11100110010111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00110001100001010000010100010011",                                                                                                
"11100101100111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00110110000001010000010100010011",                                                                                                
"11100100110111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00111010100001010000010100010011",                                                                                                
"11100100000111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"00111111000001010000010100010011",                                                                                                
"11100011010111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01000011100001010000010100010011",                                                                                                
"11100010100111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01001000000001010000010100010011",                                                                                                
"11100001110111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01001100100001010000010100010011",                                                                                                
"11100001000111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01010001000001010000010100010011",                                                                                                
"11100000010111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01001011000001010000010100010011",                                                                                                
"11011111100111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01010100110001010000010100010011",                                                                                                
"11011110110111111110000011101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01010110010001010000010100010011",                                                                                                
"11011110000111111110000011101111",                                                                                                
"00000000000100000000011110010011",                                                                                                
"11111100111101000010011000100011",                                                                                                
"11111100110001000010011110000011",                                                                                                
"00000100000001111000011001100011",                                                                                                
"11111110000001000010011000100011",                                                                                                
"00000011100000000000000001101111",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01010111000001010000010100010011",                                                                                                
"11011011110111111110000011101111",                                                                                                
"11111101110001000010010100000011",                                                                                                
"11011101000011111111000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100111101000010010000100011",                                                                                                
"11100000000111111110000011101111",                                                                                                
"00000000000001010000011110010011",                                                                                                
"11111100111101000000110110100011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"00000000000101111000011110010011",                                                                                                
"11111110111101000010011000100011",                                                                                                
"11111110110001000010011110000011",                                                                                                
"11111100110001000010011100000011",                                                                                                
"11111100111001111110001011100011",                                                                                                
"00000000000000000000010100010111",                                                                                                
"01010111000001010000010100010011",                                                                                                
"11010111110111111110000011101111",                                                                                                
"11111101110001000010010100000011",                                                                                                
"11100010010111111111000011101111",                                                                                                
"00000000000000000000011110010011",                                                                                                
"00000000000001111000010100010011",                                                                                                
"00000011110000010010000010000011",                                                                                                
"00000011100000010010010000000011",                                                                                                
"00000100000000010000000100010011",                                                                                                
"00000000000000001000000001100111",                                                                                                
"01010010010101000000110100001010",                                                                                                
"00001101000010100101000001000001",                                                                                                
"00000000000000000000000000000000",                                                                                                
"01010010010011110100001001000001",                                                                                                
"00000000000011010000101001010100",                                                                                                
"01010100010010010101100001000101",                                                                                                
"00000000000000000000110100001010",                                                                                                
"01101100011100000110110101001001",                                                                                                
"01101110011001010110110101100101",                                                                                                
"01100001011011010010000001110100",                                                                                                
"00101001001010000110111001101001",                                                                                                
"01101111011001100010000000101100",                                                                                                
"00000000000010100010000101101111",                                                                                                
"01001110010010010101101100100000",                                                                                                
"00100000010111010100111101000110",                                                                                                
"01110011011000010110110001000110",                                                                                                
"01000100010010010010000001101000",                                                                                                
"00000000000000000000000000111010",                                                                                                
"00111010011001100011000100100000",                                                                                                
"00110000001110100011011000111000",                                                                                                
"00000000000000000000000000110001",                                                                                                
"00111010011001100110001000100000",                                                                                                
"00111000001110100011010100110010",                                                                                                
"00000000000000000000000001100100",                                                                                                
"00111010011110000111100000100000",                                                                                                
"01111000001110100111100001111000",                                                                                                
"00000000000000000000000001111000",                                                                                                
"01100001011011000100011000100000",                                                                                                
"01101001001000000110100001110011",                                                                                                
"01101001011101000110100101101110",                                                                                                
"01111010011010010110110001100001",                                                                                                
"00001010001000000110010001100101",                                                                                                
"00000000000000000000000000001101",                                                                                                
"01001110010010010101101100100000",                                                                                                
"00100000010111010100111101000110",                                                                                                
"01111001011100000110111101000011",                                                                                                
"00100000011001110110111001101001",                                                                                                
"00110000001101010011001000100000",                                                                                                
"01100110001000000100001001001011",                                                                                                
"00100000011011010110111101110010",                                                                                                
"01110010011001000110010001100001",                                                                                                
"00111010011100110111001101100101",                                                                                                
"00110000011110000011000000100000",                                                                                                
"00110000001100000011000000110000",                                                                                                
"00001101000010100010111000110000",                                                                                                
"00000000000000000000000000000000",                                                                                                
"00001101000010100000110100001010",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00101101001011010010101100100000",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101011001011010010110100101101",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01000111010001010101011000100000",                                                                                                
"01100101010100110010000001000001",                                                                                                
"01110011011001010110100101110010",                                                                                                
"00100000011001100110111100100000",                                                                                                
"01110010011000110110100101001101",                                                                                                
"01101111011100100111000001101111",                                                                                                
"01110011011100110110010101100011",                                                                                                
"00100000011100110111001001101111",                                                                                                
"01100101011101100110010101000100",                                                                                                
"01100101011100000110111101101100",                                                                                                
"01111001010000100010000001100100",                                                                                                
"01000100001011010100001100100000",                                                                                                
"00100000001011000100001101000001",                                                                                                
"01001001010001000100111001001001",                                                                                                
"00100000001000000010000001000001",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"01001101001000000010000000100000",                                                                                                
"01101111011100100110001101101001",                                                                                                
"01100011011011110111001001110000",                                                                                                
"01101111011100110111001101100101",                                                                                                
"01100101010001000010000001110010",                                                                                                
"01101111011011000110010101110110",                                                                                                
"01101110011001010110110101110000",                                                                                                
"01110010010100000010000001110100",                                                                                                
"01100001011100100110011101101111",                                                                                                
"00101100011001010110110101101101",                                                                                                
"01101110011101010100011000100000",                                                                                                
"00100000011001000110010101100100",                                                                                                
"01001101001000000111100101100010",                                                                                                
"01011001011101000110100101100101",                                                                                                
"01101111010001110010000000101100",                                                                                                
"00100000001011100111010001110110",                                                                                                
"01001001001000000110011001101111",                                                                                                
"01100001011010010110010001101110",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"01000010001000000111110000100000",                                                                                                
"01101100011101000110111101101111",                                                                                                
"01100101011001000110000101101111",                                                                                                
"01110110001000000010110001110010",                                                                                                
"00110001001000000111001001100101",                                                                                                
"00110000001011100011000000101110",                                                                                                
"00100000001000000101101100100000",                                                                                                
"01100111011001000110100000101000",                                                                                                
"01100001011001000110001101000000",                                                                                                
"01110110011101000101111101100011",                                                                                                
"01010100001000000010100101101101",                                                                                                
"01001111001000000110010101110101",                                                                                                
"00100000001000000111010001100011",                                                                                                
"00110001001000000011010100110001",                                                                                                
"00110000001101010011101000110110",                                                                                                
"00100000001100100011001100111010",                                                                                                
"00100000010101000101001101001001",                                                                                                
"00110100001100100011000000110010",                                                                                                
"00110011001100010010001100100000",                                                                                                
"01111100001000000101110100110101",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"00100000010111110101111101011111",                                                                                                
"01011111001000000010000000100000",                                                                                                
"01011111010111110101111101011111",                                                                                                
"01011111010111110101111101011111",                                                                                                
"01011111010111110101111101011111",                                                                                                
"01011111010111110101111101011111",                                                                                                
"01011111010111110101111101011111",                                                                                                
"01011111010111110101111101011111",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01010011010010010010000000100000",                                                                                                
"00111010001000000010000001000001",                                                                                                
"01010011010010010101001000100000",                                                                                                
"00100000010101100010110101000011",                                                                                                
"00110011010101100101001001011011",                                                                                                
"01011101010011010100100100110010",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"01111100001000000101111101011111",                                                                                                
"00100000001011110010000000100000",                                                                                                
"00100000010111110101111100101111",                                                                                                
"01011111010111110101111100100000",                                                                                                
"00100000010111110010111101011111",                                                                                                
"01011111010111110101111100100000",                                                                                                
"01011111010111110010111101011111",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000001111100",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"01111100001000000101111101011111",                                                                                                
"00101111001000000010111100100000",                                                                                                
"00100000001000000101111101011111",                                                                                                
"00100000001011110101111101011111",                                                                                                
"00100000001000000101111100100000",                                                                                                
"01011111010111110010000000101111",                                                                                                
"00100000010111110101111100100000",                                                                                                
"00100000011111000010111100100000",                                                                                                
"00100000001000000010000001111100",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01010000010000110010000000100000",                                                                                                
"00111010001000000010000001010101",                                                                                                
"01000111010001010101011000100000",                                                                                                
"01010100010001010010000001000001",                                                                                                
"00110101001100110011000000110001",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"01111100001000000101111101011111",                                                                                                
"00100000001011110010000000101111",                                                                                                
"00101111001000000010000001011111",                                                                                                
"00100000010111110101111101011111",                                                                                                
"00101111001000000010111100100000",                                                                                                
"00101111001000000010111101011111",                                                                                                
"00100000001000000101111100100000",                                                                                                
"00100000010111110101111101011111",                                                                                                
"00100000001000000010000001111100",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"01011111010111110101111101011111",                                                                                                
"00100000001000000010111101011111",                                                                                                
"01011111010111110101111100101111",                                                                                                
"00100000001011110101111101011111",                                                                                                
"01011111010111110101110000100000",                                                                                                
"00100000001011110101111101011111",                                                                                                
"00101111010111110010111100100000",                                                                                                
"01011111011111000010000000100000",                                                                                                
"00100000001000000010000001111100",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00101101001011010010101100100000",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010101100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101101001011010010110100101101",                                                                                                
"00101011001011010010110100101101",                                                                                                
"00000000000000000000110100001010",                                                                                                
"00100000001000000111110000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01110111001000000010000000100000",                                                                                                
"01110110001011100111011101110111",                                                                                                
"01110000011000010110011101100101",                                                                                                
"01100101011000110110111101110010",                                                                                                
"01110010011011110111001101110011",                                                                                                
"01101110011010010010111001110011",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000111110000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01110110001000000010000000100000",                                                                                                
"01000000011000010110011101100101",                                                                                                
"01100011011000010110010001100011",                                                                                                
"00100000011011100110100100101110",                                                                                                
"00100000001000000010000000100000",                                                                                                
"00100000001000000010000000100000",                                                                                                
"01111100001000000010000000100000",                                                                                                
"00000000000000000000110100001010",                                                                                                
"01010100001000000000110100001010",                                                                                                
"01110011011011100110000101110010",                                                                                                
"00100000011100100110010101100110",                                                                                                
"01100101011001000110111101101101",                                                                                                
"00100000001110100000100100100000",                                                                                                
"01010100010100100100000101010101",                                                                                                
"01001111010011010101100000100000",                                                                                                
"00001010010011010100010101000100",                                                                                                
"00000000000000000010000000001101",                                                                                                
"01001001001000000000110100001010",                                                                                                
"00001001010011010100000101010010",                                                                                                
"01011011001000000011101000001001",                                                                                                
"00110000001100100111100000110000",                                                                                                
"00110000001100000011000000110000",                                                                                                
"00110000001000000010110100100000",                                                                                                
"01000110001100110011001001111000",                                                                                                
"01011101010001100100011001000110",                                                                                                
"00110101001100100101101100100000",                                                                                                
"01000010010010110010000000110110",                                                                                                
"00100000000011010000101001011101",                                                                                                
"00000000000000000000000000000000",                                                                                                
"01010000001000000000110100001010",                                                                                                
"01110011011000010110010101101100",                                                                                                
"01100101011100110010000001100101",                                                                                                
"01100110001000000110010001101110",                                                                                                
"00100000011001010110110001101001",                                                                                                
"01101110011010010111001101110101",                                                                                                
"01001101010110000010000001100111",                                                                                                
"01001101010001010100010001001111",                                                                                                
"01100100011011100110000100100000",                                                                                                
"01100101011010000111010000100000",                                                                                                
"01110010011100000010000001101110",                                                                                                
"00100000011100110111001101100101",                                                                                                
"01000101010101000100111001000101",                                                                                                
"01100101011010110010000001010010",                                                                                                
"00001101000010100010111001111001",                                                                                                
"00000000000000000000000000100000",                                                                                                
"01010011001000000000110100001010",                                                                                                
"01110100011100100110000101110100",                                                                                                
"00100000011001110110111001101001",                                                                                                
"01100111011011110111001001110000",                                                                                                
"00100000011011010110000101110010",                                                                                                
"00001010001011100010111000101110",                                                                                                
"00001010000011010000101000001101",                                                                                                
"00001010000011010000101000001101",                                                                                                
"00000000000000000000000000001101"                                                                                                                                                                                           
);
begin

	process(clk,rst_n)
	begin
		if rst_n='0' then
				
				douta <= x"00000000";     
				doutb <= x"00000000";
		
		else
			if clk'event AND clk = '1' then
			
				if  ena = '1' then
					douta		<=	CDAC_rom(conv_integer(addra(12 DOWNTO 0)));
				end if;  
				
				if  enb = '1' then
					doutb		<=	CDAC_rom(conv_integer(addrb(12 DOWNTO 0)));
				end if;
				
			end if;	
		end if;
	end process;

				            
end ROM_THEJAS32_a;          